library verilog;
use verilog.vl_types.all;
entity matarsak is
end matarsak;
